d8:announce36:http://bt1.archive.org:6969/announce13:announce-listll36:http://bt1.archive.org:6969/announceel36:http://bt2.archive.org:6969/announceee7:comment682:This content hosted at the Internet Archive at https://archive.org/details/android-x86-4.3-20130725_201512
Files may have changed, which prevents torrents from downloading correctly or completely; please check for an updated torrent at https://archive.org/download/android-x86-4.3-20130725_201512/android-x86-4.3-20130725_201512_archive.torrent
Note: retrieval usually requires a client that supports webseeding (GetRight style).
Note: many Internet Archive torrents contain a 'pad file' directory. This directory and the files within it may be erased once retrieval completes.
Note: the file android-x86-4.3-20130725_201512_meta.xml contains metadata about this torrent's contents.10:created by15:ia_make_torrent13:creation datei1654234431e4:infod11:collectionsl43:org.archive.android-x86-4.3-20130725_201512e5:filesld5:crc328:34673ab76:lengthi208666624e3:md532:8a905507c511899b109a505d8e14f2635:mtime10:14491530314:pathl28:android-x86-4.3-20130725.isoe4:sha140:b2b4ba3da4b90e9a95bfa0a088bcaa8eb5ce0c30ed5:crc328:205d61146:lengthi9216e3:md532:a3faff402bd0519370d49ec3498d9a255:mtime10:14491530494:pathl43:android-x86-4.3-20130725_201512_meta.sqlitee4:sha140:071954eb37e307145e6f1496cfbd68dd50c24a6bed5:crc328:58df48136:lengthi930e3:md532:3b34a1448c62b826b3e048223cb090c95:mtime10:16542344304:pathl40:android-x86-4.3-20130725_201512_meta.xmle4:sha140:08839f25b6de9e0d2533cc115febb3acbe8a637bee4:name31:android-x86-4.3-20130725_20151212:piece lengthi524288e6:pieces7980:�"��M�Ђ�e$g������l���U=�a��j��2`�����n4�c4k���۞�㠜�X�b��/�r�/��0��W�
�1���R�ݤvqWt��}8�p�Fg������v�̿�,�aG��_e��������I=&�ζ\Lx��|c�y�����Ͽfqu��
 :5���X��J���
����=�{CH�ld�M�.3#�)�av"v:Ů���B��Sw��TP�j��j�Y��9��1m�q�I1/>�^���tl����w��ɺX�}}��.��+��3���?":�JD��hB]q1)���M&(P��d��̳�L2Y�]�	=��n'�c<
�XT�y)���u�nЅ(V�a<�s�u�)���{������h���SU�]��^�pq��|��<@\U�$��<J����`AIp�<�����D�wO<r��䕠c9߳�1�y���On��XX��/�\�f�Y����8?N���()�	�m����n;�Z�aS�gy���K �_��MV�$|���AA-���V�C.����ʲ�,>�D��Z�W��Zq�(��ƚ������Y���Tc�ɍPF�UTE��b�J��<�9(��u��>��d���u��6�������� ��`�4&�������UU3D1�nxp���]o��ѣ���2��^[[;����l����6m�)	o��j+(�F{���h\4!��;0������l�L�vy� �� ��7����=l���`���I��E �\��.~�1����L���=�+꾦Kk;hQ�������W�+�<���.ͧ_�~b��|����N��fՅ�i�0��o�p�F��Y�cι��	m����sg{�jX��l�%q$g�t�w3���[�2�����|� ���r ֽ����N}/�=�vnd ��WQVX�U���;3�@F4�vⶌ������_c(���b��ׇ���P_�d�����b7���_+G��M�eU-��oN�~�|�V���T�����Μ�O�V�>�D��hO2��sf~�J�d+��1y��;��+�N�K���O^����0õ;4yZ-�GG^x��=����9P�^������X��Tx-/y0�Rj�u(���N���g�;e�SIGb�h�����C��3!@��p����bU+��߻q��a���[�k��jM�ƆS�����{_��S��+�^��s�)����n6�tܗ�4-ޚ'�c��d�'��WK,���=ӝ��$�6dP?�l�X��'�:��ҝ���I��Z����)�M�q��(�'<a�1����W�W�H{)dQ<HA��GH��ܡ:ϭ\�sG+��mv��&�E�lD6$�Db�L�q#�Ӹy�3���4(�r�20b�ȝAO�7��)r|��-���Q�-jR�s&M�|����0��� �5���O�Ȕ׈E�`*��|/7>�BȣLu��"���	����k�E�6�S�5Š�	v@b~2�,����rhP��Uz)��x�� Q�B;?���W��_)�v<�9Zݨy�DǇ�jEF?l��pe����w�����>�:dik\3I	��@|m	x03gh��6=�TW��ɤV=��o�QASV:7c�7陳�+I~�x�7]������@����9����!P�_�:3��"x���cPo��.�O���4Y3<cY�<g��� ���Va�ʟ��x��	��zN�$v��B�K��@Q^�n�[�K�߄X�+Ir�Mmm���[����׭���D�� ����р��6QjpG�~�pP�<������o�|ߡ���ϟr1�6�	Tqv��ܗ����x���*UQ�����s���_]�竛^�Ck�4;�U����=�ӚE�)����*N�4����9��p.aq��.�v���m=�����Ρζ�d�������k��h���X�0O�c����{:��<��jF>\C��|�V5J$�`Thi�EO��a*�j����gU���ӷ� /�Wytxɩ��	�{����,�l�-�~�*Y�T
\wN��	�8AX�;Z`6����4�g�|Ė�M�ۛڠ�v�+ė
ݷ��N�z]{��>�|$��Lӿ1�P<ڠD�Z����/���g7o���Z��5)�H�[=!�z�B���\f���?o��n@���\c�o3O�7��� E<[�8�,���4��]Y�\�`�N픍)ɻC�J�&4n_��6ԐF�{tC'��<�h���A,�Iu�w5��n2Ԓ^���1�K�����~'�D�G�����	H� 7FD(t���^�_cOג���J���-bO&�'$�����6H��<^_4�QU�w�F�}�%w=���BZÔ�L��/�T��>�^ڒ���
$s|�4Q64兎� �Qa+&m�:xDtiPe%A̭�~J�k�T�	�ڔ"����X���߁�ݳ4ެў	�I~4&v3� �{¦moc¦;U�AqJ�h-�>�M�e8��;�X�(%�/_БG���y�?G!`i���c`,ax�F4-�7�
�xj}"�����Ã5�˻�k�[�+���g����g�81z�ύ�^_3�4��9��s%o~��)~u�_-�����m�i�z����52	���=4|Z#c��MeM����t��_���Fؔ� ��XDq|F=̙?\��顥(�T�$K2~�YSy����e�W�T:�="כI�~�ڈ�p��E���R��Ǎ/<i��OӐ�;���^����J���V#�� 2�%�3$�e�=�p�*�?�s겯ĥ�J��Td�7��XK!S�[�H�>���K6{�Or.��`|��B(�(�;\�x��D��<Ak;Y�ރu��/S):xqi��N�%*$Ҭ���:�g��걠!O�9��L�
��Y��9���f�2yvW�΢�����u��%b[�3�:	ˋS�4�1��xs�O������>�[��T��6u���`�������
9�oX.��4�?��y�;�	�����k���tX#0EҮ�b���:>���C&=[ٺ���a�#4��$
	�����B��6��ĸ���e�x��˗�����2_�xQ�������ۿ������\4���H§a!�_Ú�Q�[2m���ٲ �0[*��V�m���ݑ�&�R;}�Ϋ�*D��G W��%���N��.�ҦK��|<̔�Me��H��}J�$�^a]�������K�	v�Ù&�뿿:1���2!"C�3PQ-�s�'TD=����eK�셙��l2��oI��S����;gF%F/PdR!W��R0Y� QS�]���7zs�E��$߾���?���ϩ�� ���� ����	߹U�3�o�Εx`��
�a��'ߐ���.��`TS�����_�ߢ� x�W�����=f�ٟԌz`�Z�%��{��!
U�Ml��)ᏼ�< Lڜ��&_8X�K.2���H�u�!��Sc��2;��;O����c�|�o!Ok�Y%x҂^x��fk]�<��_���L����x6Y5p��x��ü�}7�[$v�0{8�8�t!(76#I͏^<3�0C�����?�֍�����W�|�>�;� ih��CSA7�^x?_��������n��u��β�m�#�����	���󑖶:�	���r�a��N	��F#�n&?�mbL���`�y�l��3���=zofOꐇ�g� 0h`���$&�_nj�%���_Y d6���Z��kw��p���=$b�i��[��"�^۽qh�>@�>�w�^�^٦7BO	�?���hr��p��c�
���{QAk4{�C&�`���Y�^�\� \9heGr�ŭ޷҉i�d�ߣH�2֨n5q�D��#��(^�m�J,p�Wp�'�wԓ����I��<)�SLP�^qD�rjA4:L�&J�s/#&�L�f`�;��0�@���:�/ڬ^���)��ѷ$Z�0dQ���g=�2��~J9��kk�l���|������m�1�'�v��>�P��m��u09^�@�,5�on?�`S����齷Ҽ�J^�V��L�1��r^ �V\mn����w���p�A��*��h�X��3��	a�>�"_c|�-��ض46�p����W7g�A���W���y��?ߕ��?o&L��#zb�펣y�͊"��O�e��yP+�[<nK���v"�W�ޖ��^{�j�Ey���#��EcU�y	�&~�^Y�7�J�&���&���\q�ցs�y
s�V�Iaq�C$"�Bp���� ��?>E���c#mѬ	f~ݤ�Jr�]x��:,h�r��2�]���}J*W%w�te�+��U��v7�����J�M�P��|�U@?�b&��!m��Vu�F)��L8���K�(Y��@�i�� �Z�֒:��P#.E��.} >�@I��5=]�KR�'6[Aو��.���Ʌʅ���8�G ��2mZ��E�n׆h�u��$���v2B��d���5m�N�4�z��)I@�}D�L��+��kkx�$�x�Ț�Z#�?���e�kɇ�6��>�xx�(b��U1@Y)z�?�c�y�U����9�,����F'/ã7�VE�FoY� <��i�a��pUL�x�u�mK�?��ⲔÎϪu�Op�D�x�{T�Iܖ}�(�5N|C	�?\ӭX�����x�x�i�j�+��N�����#{�a�ǃi��E. �-�F%�1z�Tk�mBME���-]9잧�c�<����5�@8ގ:=�Q�����'0��l��B�[���f�ҩ��MǇ��?y�=��t�f��G7����SU��iåQ����9�٫$�f8��o�VPU�g��m�	��־� ��%\�;}�Ų9[�{�z�v[��	=_��Y���J��W�s����)8�~r�-��aA���bq E�%$&��E��$m�"���$�XlS<�ڭd�ZX�%O2iƄ�z
�0-��rʚ��+�Z���^����O�'�D	@�x.���)����	�!;�)!:U� ְ�� Un ��D�k�"M���Ra�������w1Ⱦ�H��V���i����,i�/G��K�j�7��N-IQ��؍�:ܒ�ҭ�?G3�:�� Ì��e\������I��˼,/c�j�#�l���ĥs��M�Ζ���/�����ܗ�Xi;U�K���|�ު_�����QG^]+c��A6�.]�we�쐾�B��TK�C�G}";�| H�ص�Id�#�5�f����@�� �'f�԰� |>�9�_]�����1��8X]k��.���gE}��ڳ����ӈ�Bu]\���FŊʽˇ�`���u�J��jD���oķEQ�P>f�}�$�ђ�fk�Ӷ�=IL*h�����lꛑ>�da�<�dYl����pBX�Brrױ)u8'�t����gCK�QqF��{>�03��O���O�dD6ӝ��'�7M7�9j��J'#D,�Ziw�g`P5x�&K�9��ģ,�Y����2q����0!.���[;dW~�%7���6u ���i�{�R]A��b䉝����]Z�������;���u�k��tYW�c�1���5�L6H�̢ q�LZW�u��q��}gu�U,.խ��~�쩐�[X��`��dɝbL�5*S7V�#�"���yِ4���5�Xs��ө�9H��HS<��AM���Q��<�Ӥ�ɅxU���*���( �+������9��H��*��$�D�%9�!F e�<*Jr!��%�å@�c�<����51��"�T��Zy�+�j*4���C���o�c���O�,�e\!�#��6��
���(>�䌴��)�=.�#�B��Ǿ1�]\!�TM�T� ��tyT��]h�ҟk���Ũc�rmu1�N5�WI��\�-���`�m3�z6�[Z'�adW�0�7��H:F�r�����v����Ggxk��\ȧK��E�ח��6����A��i[��F����o���t:�kj=
]Q��zaG��J�Z3�&�Ό���ML��D��^E�̿2v���)���0�Ҽ3im1�������J;�x�o6˼e�
1Xk����yI���3k��a�������t�YSB�q�\�[�p����%�;�mn�=��4y;��x@͌�G���� �#��2���ONtMPGK���;%�R�,����s�@0!����bzNK���̆ ���9���Gї�Gq|�c��]_�0� ��W������R+̿��j��&�����i	494$q^/�dvF�^�%�$�f{x��``���M�E��ap��-Lg}���_ʽ]K���V�&�/Eϑ4�m��3G�Y(T�!o�� NS�D�&�A���R��L6͉�p���쀩�ab�i�"�ul;��� 
騥�������� HQx��"X�V�K�l����_\y	�盷����v��<Ⱦ�	�ok�=�pu����q�)�T*�����ܬ�5��OI�՛�c����n���Cy�J.9�
ۣh&8O$,���~]�:�-�'H�'>�ڞI=/4��S�6*�e����G�
�m�l	��<��4������Ņcq�cڹ��!C�y����]xI�N��|����C�����]�ߐC
]��-8����d;�O"'�Qpg�y)��4)@������:d6��jS˖U�Fj�y�ݻJL
'�%�0҄N���ĻK�T��A�0���@ԙ �X��!�|��X!o�ӗ��`@���7�qCy�53���g�6�N����wc�ye�[��Z�]��������*e���'t'<�5G�gyGl����?�i��@](�+\z�9����^��!����bipP���
��=NɃ!����ՕO��\�p
�����7�Į�??�$�o���X�GA�V^"���+,}A�ws�h��~��urxLT�=���=�#�*O-^�:(��xI���m���Tyo?�h�����B��ϾU�Bw�S`�Y�/j��Y��tE��$`^�F�<8��y��;�cS���Y�տvkg-P��L�Bˑ�c�-,��ȼ`�Y��a҆N��r���R)*��� \�|����Yf��i>�<���l0,~@y����FJj�)I%�l�����E;�xo�5ξ�Kο_��]�GZQ,'A&:7���ߵ;5��.vg���*�&i�L�
&�����}Z��ݬ��I"v��Z�m����%�+�02/�BB|�q������K���l2N�+���d�cs#C��neI ��^�s�=���<��i�]W��ˌ�w*�<8�s��F��,% @���h�A�@Xg��v�Ԩ9����nz{m���c+�A_�_J�0���!FТf�=��cԘ�Z�5噻ȱP��k��`��'3&�b�RD�x~�,��0�������i�,�PXU ��`	�؋��X��f�l`U"UG 	���nb��bϱWtY����ļ���W4�Ŷ�]ߤ�WT:)z��n�뒉6�_EŒ<��3G]Ĥ�P8���'$hު�����c(M�x[i��`�?�yv0�)H�<}m����BJi��Ln\r�{�v�e6��|n�K�����ad��%�
i���(9���2p:�T�q���N��_A���O/�'��
P�;3ȼx�/��L��}]b�vyC��vq>�:��uYdQI
R�m�+��ǋ�o�-�&b7��Cʗ�"���J"�-d�J[�w`�C�F.�?�4?����f�p�)�-`ê����^ 9�V�Ho�*:�(嬺s������^8ޢ�R+6��/�q=��P/�P��5Z�WjR*c,&�;���K���挘ڏ��N����y�i�Y-e6:locale2:en5:title31:android-x86-4.3-20130725_2015128:url-listl29:https://archive.org/download/40:http://ia601304.us.archive.org/16/items/10:/16/items/ee